module Nand_Gate(out,in1,in2);
  
  input in1,in2;
  output out;
  
  nand(out,in1,in2);
  
endmodule
