module Not_Gate(out,in);
  
  input in;
  output out;
  
  assign out = !in;
  
endmodule