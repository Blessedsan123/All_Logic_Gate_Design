module Nor_Gate(out,in1,in2);
  
  input in1,in2;
  output out;
  
  nor(out,in1,in2);
  
endmodule