module Xor_Gate(out,in1,in2);
  
  input in1,in2;
  output out;
  
  xor(out,in1,in2);
  
endmodule