module Xnor_Gate(out,in1,in2);
  
  input in1,in2;
  output out;
  
  xnor(out,in1,in2);
  
endmodule